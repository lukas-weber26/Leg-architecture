module LEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_15), .en(wire_48), .out(arch_output_value));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_1 (.en(wire_33), .in(arch_input_value), .out(wire_28));
  TC_Or # (.UUID(64'd3157105682597732050 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_56), .in1(wire_5), .out(wire_64));
  TC_Or # (.UUID(64'd700045591590561234 ^ UUID), .BIT_WIDTH(64'd1)) Or_3 (.in0(wire_58), .in1(wire_27), .out(wire_115));
  TC_Or # (.UUID(64'd3549001667251634900 ^ UUID), .BIT_WIDTH(64'd1)) Or_4 (.in0(wire_50), .in1(wire_19), .out(wire_66));
  TC_Or # (.UUID(64'd2269694454788292946 ^ UUID), .BIT_WIDTH(64'd1)) Or_5 (.in0(wire_74), .in1(wire_14), .out(wire_86));
  TC_Or # (.UUID(64'd1844048388294245364 ^ UUID), .BIT_WIDTH(64'd1)) Or_6 (.in0(wire_62), .in1(wire_45), .out(wire_101));
  TC_Or # (.UUID(64'd2695359556586327911 ^ UUID), .BIT_WIDTH(64'd1)) Or_7 (.in0(wire_67), .in1(wire_34), .out(wire_113));
  TC_Switch # (.UUID(64'd2646728809043152279 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_56), .in(wire_40), .out(wire_17_0));
  TC_Switch # (.UUID(64'd1935160467439464196 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_5), .in(wire_40), .out(wire_2_8));
  TC_Switch # (.UUID(64'd977321102049953818 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_58), .in(wire_106), .out(wire_17_2));
  TC_Switch # (.UUID(64'd3722515247921723471 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_27), .in(wire_106), .out(wire_2_7));
  TC_Switch # (.UUID(64'd3601188592565593964 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_50), .in(wire_97), .out(wire_17_4));
  TC_Switch # (.UUID(64'd4014399076376933194 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_19), .in(wire_97), .out(wire_2_6));
  TC_Switch # (.UUID(64'd4161672925644182449 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_74), .in(wire_73), .out(wire_17_3));
  TC_Switch # (.UUID(64'd552375585198440410 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_14), .in(wire_73), .out(wire_2_5));
  TC_Switch # (.UUID(64'd4265176839667625262 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_62), .in(wire_79), .out(wire_17_5));
  TC_Switch # (.UUID(64'd1041730340393858558 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_45), .in(wire_79), .out(wire_2_4));
  TC_Switch # (.UUID(64'd491192510242440390 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_67), .in(wire_32), .out(wire_17_6));
  TC_Switch # (.UUID(64'd2442295756390004600 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_34), .in(wire_32), .out(wire_2_1));
  TC_Or # (.UUID(64'd4129098185517505965 ^ UUID), .BIT_WIDTH(64'd1)) Or_20 (.in0(wire_71), .in1(wire_42), .out(wire_33));
  TC_Switch # (.UUID(64'd2312725337422069148 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_71), .in(wire_28), .out(wire_17_8));
  TC_Switch # (.UUID(64'd3907588151097613508 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_42), .in(wire_28), .out(wire_2_2));
  TC_Switch # (.UUID(64'd2410113394107929429 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_83), .in(wire_9), .out(wire_17_7));
  TC_Switch # (.UUID(64'd1826964660860977844 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_75), .in(wire_9), .out(wire_2_0));
  TC_Add # (.UUID(64'd1836364419457964329 ^ UUID), .BIT_WIDTH(64'd8)) Add8_25 (.in0(wire_1), .in1(wire_13), .ci(1'd0), .out(wire_69), .co());
  TC_Decoder3 # (.UUID(64'd4598855726905540096 ^ UUID)) Decoder3_26 (.dis(wire_91), .sel0(wire_54), .sel1(wire_120), .sel2(wire_104), .out0(wire_56), .out1(wire_58), .out2(wire_50), .out3(wire_74), .out4(wire_62), .out5(wire_67), .out6(wire_83), .out7(wire_71));
  TC_Decoder3 # (.UUID(64'd388667379281544807 ^ UUID)) Decoder3_27 (.dis(wire_90), .sel0(wire_124), .sel1(wire_100), .sel2(wire_135), .out0(wire_5), .out1(wire_27), .out2(wire_19), .out3(wire_14), .out4(wire_45), .out5(wire_34), .out6(wire_75), .out7(wire_42));
  TC_Decoder3 # (.UUID(64'd1926417040054614309 ^ UUID)) Decoder3_28 (.dis(wire_122), .sel0(wire_127), .sel1(wire_80), .sel2(wire_96), .out0(wire_8), .out1(wire_35), .out2(wire_51), .out3(wire_29), .out4(wire_110), .out5(wire_53), .out6(wire_37), .out7(wire_48));
  TC_Add # (.UUID(64'd918325968594195230 ^ UUID), .BIT_WIDTH(64'd8)) Add8_29 (.in0(wire_1), .in1(wire_131), .ci(1'd0), .out(wire_95), .co());
  TC_Neg # (.UUID(64'd878407423054571151 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_30 (.in(wire_13), .out(wire_131));
  TC_And # (.UUID(64'd4274290278184732434 ^ UUID), .BIT_WIDTH(64'd8)) And8_31 (.in0(wire_1), .in1(wire_13), .out(wire_16));
  TC_Or # (.UUID(64'd1547202834476000431 ^ UUID), .BIT_WIDTH(64'd8)) Or8_32 (.in0(wire_1), .in1(wire_13), .out(wire_81));
  TC_Xor # (.UUID(64'd4239535398454787880 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_33 (.in0(wire_1), .in1(wire_13), .out(wire_128));
  TC_Decoder3 # (.UUID(64'd389698951624136615 ^ UUID)) Decoder3_34 (.dis(1'd0), .sel0(wire_57), .sel1(wire_22), .sel2(wire_20), .out0(wire_25), .out1(wire_70), .out2(wire_31), .out3(wire_65), .out4(wire_52), .out5(wire_44), .out6(wire_89), .out7(wire_121));
  TC_Splitter8 # (.UUID(64'd3268803031893760400 ^ UUID)) Splitter8_35 (.in(wire_94[7:0]), .out0(wire_57), .out1(wire_22), .out2(wire_20), .out3(), .out4(), .out5(wire_77), .out6(wire_108), .out7(wire_105));
  TC_Switch # (.UUID(64'd854224910746831379 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_129), .in(wire_69), .out(wire_4_7));
  TC_Switch # (.UUID(64'd1134581407703562038 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_37 (.en(wire_117), .in(wire_95), .out(wire_4_6));
  TC_Switch # (.UUID(64'd339522117565355418 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_133), .in(wire_16), .out(wire_4_4));
  TC_Switch # (.UUID(64'd696553676050962115 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_39 (.en(wire_116), .in(wire_81), .out(wire_4_2));
  TC_Switch # (.UUID(64'd1297438585075373775 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_40 (.en(wire_99), .in(wire_128), .out(wire_4_5));
  TC_Counter # (.UUID(64'd4565566535796709893 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_41 (.clk(clk), .rst(rst), .save(wire_43), .in(wire_15), .out(wire_9));
  TC_Constant # (.UUID(64'd2421151058344302069 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_42 (.out(wire_46));
  TC_Switch # (.UUID(64'd2530858208274395553 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_43 (.en(wire_68[0:0]), .in(wire_46), .out(wire_43));
  TC_Splitter8 # (.UUID(64'd1709856727448948382 ^ UUID)) Splitter8_44 (.in(wire_21), .out0(wire_127), .out1(wire_80), .out2(wire_96), .out3(wire_39), .out4(wire_23), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd806974381889649167 ^ UUID)) Splitter8_45 (.in(wire_55[7:0]), .out0(wire_124), .out1(wire_100), .out2(wire_135), .out3(wire_6), .out4(wire_10), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd2700067647918424519 ^ UUID)) Splitter8_46 (.in(wire_0[7:0]), .out0(wire_54), .out1(wire_120), .out2(wire_104), .out3(wire_12), .out4(wire_24), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3033746027149519320 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_85), .in(wire_17), .out(wire_1_0));
  TC_Switch # (.UUID(64'd4294820733219689153 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_119), .in(wire_0[7:0]), .out(wire_1_1));
  TC_Not # (.UUID(64'd1597131477542014239 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_105), .out(wire_85));
  TC_Switch # (.UUID(64'd3052144910283265517 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_125), .in(wire_2), .out(wire_13_1));
  TC_Switch # (.UUID(64'd1741968484046812876 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_108), .in(wire_55[7:0]), .out(wire_13_0));
  TC_Not # (.UUID(64'd1831175443725239523 ^ UUID), .BIT_WIDTH(64'd1)) Not_52 (.in(wire_108), .out(wire_125));
  TC_Not # (.UUID(64'd1041162876508567575 ^ UUID), .BIT_WIDTH(64'd1)) Not_53 (.in(wire_85), .out(wire_119));
  TC_And # (.UUID(64'd2870657483632612144 ^ UUID), .BIT_WIDTH(64'd1)) And_54 (.in0(wire_36), .in1(wire_25), .out(wire_129));
  TC_Not # (.UUID(64'd1051407927069804865 ^ UUID), .BIT_WIDTH(64'd1)) Not_55 (.in(wire_77), .out(wire_36));
  TC_And # (.UUID(64'd2760458169754153360 ^ UUID), .BIT_WIDTH(64'd1)) And_56 (.in0(wire_36), .in1(wire_70), .out(wire_117));
  TC_And # (.UUID(64'd401520817493034818 ^ UUID), .BIT_WIDTH(64'd1)) And_57 (.in0(wire_36), .in1(wire_31), .out(wire_133));
  TC_And # (.UUID(64'd498821885646581480 ^ UUID), .BIT_WIDTH(64'd1)) And_58 (.in0(wire_36), .in1(wire_65), .out(wire_116));
  TC_And # (.UUID(64'd2447005432645015302 ^ UUID), .BIT_WIDTH(64'd1)) And_59 (.in0(wire_36), .in1(wire_44), .out(wire_99));
  TC_Equal # (.UUID(64'd2595345319306895954 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_60 (.in0(wire_1), .in1(wire_13), .out(wire_82));
  TC_Equal # (.UUID(64'd3703368834552926204 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_61 (.in0(wire_1), .in1(wire_13), .out(wire_63));
  TC_Not # (.UUID(64'd444900149187627701 ^ UUID), .BIT_WIDTH(64'd1)) Not_62 (.in(wire_63), .out(wire_114));
  TC_LessU # (.UUID(64'd846358567681372337 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_63 (.in0(wire_1), .in1(wire_13), .out(wire_130));
  TC_LessU # (.UUID(64'd4378439148176752740 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_64 (.in0(wire_1), .in1(wire_13), .out(wire_107));
  TC_Or # (.UUID(64'd2571598757259102472 ^ UUID), .BIT_WIDTH(64'd1)) Or_65 (.in0(wire_107), .in1(wire_41), .out(wire_103));
  TC_Equal # (.UUID(64'd414073839477721741 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_66 (.in0(wire_1), .in1(wire_13), .out(wire_41));
  TC_Not # (.UUID(64'd2596639727405805731 ^ UUID), .BIT_WIDTH(64'd1)) Not_67 (.in(wire_26), .out(wire_88));
  TC_LessU # (.UUID(64'd519372185152537649 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_68 (.in0(wire_1), .in1(wire_13), .out(wire_87));
  TC_Not # (.UUID(64'd2248732738014538350 ^ UUID), .BIT_WIDTH(64'd1)) Not_69 (.in(wire_87), .out(wire_78));
  TC_LessU # (.UUID(64'd1604112865851423542 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_70 (.in0(wire_1), .in1(wire_13), .out(wire_26));
  TC_And # (.UUID(64'd3945878599032359685 ^ UUID), .BIT_WIDTH(64'd1)) And_71 (.in0(wire_88), .in1(wire_111), .out(wire_109));
  TC_Not # (.UUID(64'd4573437367456573398 ^ UUID), .BIT_WIDTH(64'd1)) Not_72 (.in(wire_132), .out(wire_111));
  TC_Equal # (.UUID(64'd2716325810528261246 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_73 (.in0(wire_1), .in1(wire_13), .out(wire_132));
  TC_Switch # (.UUID(64'd673946438953339171 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_74 (.en(wire_7), .in(wire_82), .out(wire_38_1));
  TC_Switch # (.UUID(64'd3371584292052594049 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_75 (.en(wire_47), .in(wire_114), .out(wire_38_0));
  TC_Switch # (.UUID(64'd1378792336298015330 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_76 (.en(wire_61), .in(wire_130), .out(wire_38_2));
  TC_Switch # (.UUID(64'd947531997621985833 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_77 (.en(wire_92), .in(wire_103), .out(wire_38_3));
  TC_Switch # (.UUID(64'd265481021936700343 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_78 (.en(wire_112), .in(wire_109), .out(wire_38_4));
  TC_Switch # (.UUID(64'd1971708582949430590 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_79 (.en(wire_98), .in(wire_78), .out(wire_38_5));
  TC_And # (.UUID(64'd3236879926515392645 ^ UUID), .BIT_WIDTH(64'd1)) And_80 (.in0(wire_11), .in1(wire_25), .out(wire_7));
  TC_And # (.UUID(64'd2773225214563595961 ^ UUID), .BIT_WIDTH(64'd1)) And_81 (.in0(wire_11), .in1(wire_70), .out(wire_47));
  TC_And # (.UUID(64'd4190607731312021098 ^ UUID), .BIT_WIDTH(64'd1)) And_82 (.in0(wire_11), .in1(wire_31), .out(wire_61));
  TC_And # (.UUID(64'd1448656918940484375 ^ UUID), .BIT_WIDTH(64'd1)) And_83 (.in0(wire_11), .in1(wire_65), .out(wire_92));
  TC_And # (.UUID(64'd3039291406258388458 ^ UUID), .BIT_WIDTH(64'd1)) And_84 (.in0(wire_11), .in1(wire_52), .out(wire_112));
  TC_And # (.UUID(64'd3350066253842505889 ^ UUID), .BIT_WIDTH(64'd1)) And_85 (.in0(wire_11), .in1(wire_44), .out(wire_98));
  TC_Not # (.UUID(64'd3727845057996746069 ^ UUID), .BIT_WIDTH(64'd1)) Not_86 (.in(wire_36), .out(wire_11));
  TC_Switch # (.UUID(64'd799678726905260767 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_87 (.en(wire_60), .in(wire_4), .out(wire_15_1));
  TC_Not # (.UUID(64'd4586230999365729696 ^ UUID), .BIT_WIDTH(64'd1)) Not_88 (.in(wire_11), .out(wire_60));
  TC_Switch # (.UUID(64'd3445840660294330351 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_89 (.en(wire_11), .in(wire_18[7:0]), .out(wire_15_0));
  TC_Constant # (.UUID(64'd4399458456191339621 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_90 (.out(wire_118));
  TC_Switch # (.UUID(64'd3005342052167319338 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_91 (.en(wire_11), .in(wire_118), .out(wire_21_1));
  TC_Switch # (.UUID(64'd4290267753472666013 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_92 (.en(wire_134), .in(wire_18[7:0]), .out(wire_21_0));
  TC_Not # (.UUID(64'd3825911746791069795 ^ UUID), .BIT_WIDTH(64'd1)) Not_93 (.in(wire_11), .out(wire_134));
  TC_Switch # (.UUID(64'd1715020736529367778 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_94 (.en(wire_38), .in({{7{1'b0}}, wire_37 }), .out(wire_68));
  TC_And # (.UUID(64'd1891321579910097234 ^ UUID), .BIT_WIDTH(64'd1)) And_95 (.in0(wire_36), .in1(wire_52), .out(wire_84));
  TC_Switch # (.UUID(64'd1417563971881493595 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_96 (.en(wire_84), .in(wire_126), .out(wire_4_1));
  TC_Not # (.UUID(64'd2695720571148029808 ^ UUID), .BIT_WIDTH(64'd8)) Not8_97 (.in(wire_1), .out(wire_126));
  TC_Shr # (.UUID(64'd3927377563627395232 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_98 (.in(wire_1), .shift(wire_13), .out(wire_49));
  TC_Shl # (.UUID(64'd3399905466696027778 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_99 (.in(wire_1), .shift(wire_13), .out(wire_30));
  TC_And # (.UUID(64'd1376211004588932381 ^ UUID), .BIT_WIDTH(64'd1)) And_100 (.in0(wire_36), .in1(wire_89), .out(wire_102));
  TC_Switch # (.UUID(64'd1131807739917282845 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_101 (.en(wire_102), .in(wire_49), .out(wire_4_3));
  TC_And # (.UUID(64'd741833455100237819 ^ UUID), .BIT_WIDTH(64'd1)) And_102 (.in0(wire_36), .in1(wire_121), .out(wire_93));
  TC_Switch # (.UUID(64'd4536640796151389046 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_103 (.en(wire_93), .in(wire_30), .out(wire_4_0));
  TC_Switch # (.UUID(64'd1628247066521983035 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_104 (.en(wire_12), .in(wire_123[7:0]), .out(wire_17_9));
  TC_Switch # (.UUID(64'd3862761475475355545 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_105 (.en(wire_6), .in(wire_123[7:0]), .out(wire_2_3));
  TC_Or # (.UUID(64'd871131906096684078 ^ UUID), .BIT_WIDTH(64'd1)) Or_106 (.in0(wire_12), .in1(wire_6), .out(wire_59));
  TC_Program # (.UUID(64'd4465777506522231470 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_3DF9A0FB422FF2AE.w8.bin"), .ARG_SIG("Program_3DF9A0FB422FF2AE=%s")) Program_107 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_9 }), .out0(wire_94), .out1(wire_0), .out2(wire_55), .out3(wire_18));
  TC_Or # (.UUID(64'd4142766655636487847 ^ UUID), .BIT_WIDTH(64'd1)) Or_108 (.in0(wire_23), .in1(wire_39), .out(wire_122));
  TC_Or # (.UUID(64'd2667232978288855861 ^ UUID), .BIT_WIDTH(64'd1)) Or_109 (.in0(wire_10), .in1(wire_6), .out(wire_90));
  TC_Or # (.UUID(64'd440214736546703614 ^ UUID), .BIT_WIDTH(64'd1)) Or_110 (.in0(wire_24), .in1(wire_12), .out(wire_91));
  TC_Switch # (.UUID(64'd3671466828535083198 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_111 (.en(wire_10), .in(wire_3), .out(wire_2_9));
  TC_Switch # (.UUID(64'd1082142112497736599 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_112 (.en(wire_24), .in(wire_3), .out(wire_17_1));
  TC_Or # (.UUID(64'd4345493239101073947 ^ UUID), .BIT_WIDTH(64'd1)) Or_113 (.in0(wire_24), .in1(wire_10), .out(wire_76));
  TC_Ram # (.UUID(64'd1193065637140015650 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_114 (.clk(clk), .rst(rst), .load(wire_59), .save(wire_39), .address({{24{1'b0}}, wire_72 }), .in0({{56{1'b0}}, wire_15 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_123), .out1(), .out2(), .out3());
  RegisterPlus # (.UUID(64'd3045777980693743268 ^ UUID)) RegisterPlus_115 (.clk(clk), .rst(rst), .Load(wire_64), .Save_value(wire_15), .Save(wire_8), .Always_output(), .Output(wire_40));
  RegisterPlus # (.UUID(64'd1157312672670656225 ^ UUID)) RegisterPlus_116 (.clk(clk), .rst(rst), .Load(wire_115), .Save_value(wire_15), .Save(wire_35), .Always_output(), .Output(wire_106));
  RegisterPlus # (.UUID(64'd263652518613353595 ^ UUID)) RegisterPlus_117 (.clk(clk), .rst(rst), .Load(wire_66), .Save_value(wire_15), .Save(wire_51), .Always_output(), .Output(wire_97));
  RegisterPlus # (.UUID(64'd2306915739580997297 ^ UUID)) RegisterPlus_118 (.clk(clk), .rst(rst), .Load(wire_86), .Save_value(wire_15), .Save(wire_29), .Always_output(), .Output(wire_73));
  RegisterPlus # (.UUID(64'd1473024321561741166 ^ UUID)) RegisterPlus_119 (.clk(clk), .rst(rst), .Load(wire_101), .Save_value(wire_15), .Save(wire_110), .Always_output(), .Output(wire_79));
  RegisterPlus # (.UUID(64'd602464059498925265 ^ UUID)) RegisterPlus_120 (.clk(clk), .rst(rst), .Load(wire_113), .Save_value(wire_15), .Save(wire_53), .Always_output(wire_72), .Output(wire_32));
  STACK # (.UUID(64'd4532388211661779513 ^ UUID)) STACK_121 (.clk(clk), .rst(rst), .POP(wire_76), .PUSH(wire_23), .VALUE(wire_15), .OUTPUT(wire_3));
  TC_LessI # (.UUID(64'd2406372620020937389 ^ UUID), .BIT_WIDTH(64'd16)) LessI16_122 (.in0(16'd0), .in1(16'd0), .out());

  wire [63:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  wire [7:0] wire_2_6;
  wire [7:0] wire_2_7;
  wire [7:0] wire_2_8;
  wire [7:0] wire_2_9;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8|wire_2_9;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_4_0;
  wire [7:0] wire_4_1;
  wire [7:0] wire_4_2;
  wire [7:0] wire_4_3;
  wire [7:0] wire_4_4;
  wire [7:0] wire_4_5;
  wire [7:0] wire_4_6;
  wire [7:0] wire_4_7;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5|wire_4_6|wire_4_7;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_13_0;
  wire [7:0] wire_13_1;
  assign wire_13 = wire_13_0|wire_13_1;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_15_0;
  wire [7:0] wire_15_1;
  assign wire_15 = wire_15_0|wire_15_1;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_17_0;
  wire [7:0] wire_17_1;
  wire [7:0] wire_17_2;
  wire [7:0] wire_17_3;
  wire [7:0] wire_17_4;
  wire [7:0] wire_17_5;
  wire [7:0] wire_17_6;
  wire [7:0] wire_17_7;
  wire [7:0] wire_17_8;
  wire [7:0] wire_17_9;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2|wire_17_3|wire_17_4|wire_17_5|wire_17_6|wire_17_7|wire_17_8|wire_17_9;
  wire [63:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [7:0] wire_21_0;
  wire [7:0] wire_21_1;
  assign wire_21 = wire_21_0|wire_21_1;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [0:0] wire_33;
  assign arch_input_enable = wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_38_0;
  wire [0:0] wire_38_1;
  wire [0:0] wire_38_2;
  wire [0:0] wire_38_3;
  wire [0:0] wire_38_4;
  wire [0:0] wire_38_5;
  assign wire_38 = wire_38_0|wire_38_1|wire_38_2|wire_38_3|wire_38_4|wire_38_5;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  assign arch_output_enable = wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [63:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [7:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [63:0] wire_94;
  wire [7:0] wire_95;
  wire [0:0] wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [7:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [7:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [0:0] wire_122;
  wire [63:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [7:0] wire_126;
  wire [0:0] wire_127;
  wire [7:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [7:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [0:0] wire_135;

endmodule
